module top(
    input clk,
    input resetn,
    axi4_Lite.axiSlave axiS_Top,
    apb.masterAPB apbM_Top
);
    converter converter(clk, resetn, axiS_Top.axiSlave,apbM_Top.masterAPB);
endmodule