module controller(
);
    
endmodule

// если в APB setup, то мы не передаем новые данные