package respone_pkg;

parameter OKAY = 2'b00; //use
parameter EXOKAY = 2'b01;
parameter SLVERR = 2'b10;   //use
parameter DECERR = 2'b11;

endpackage